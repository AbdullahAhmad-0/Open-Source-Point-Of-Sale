Demo:210.297.mm